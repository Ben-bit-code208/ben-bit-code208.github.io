#include system
module test
  import system

  func main()
	print("Hello, World!")
  end
end